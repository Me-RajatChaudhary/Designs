module SequenceDetector
