module factorial
  
endmodule
